
-- 
-- Definition of  video_buf
-- 
--      09/20/12 14:44:19
--      
--      Precision RTL Synthesis, 2012a.10
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.all;
-- Library use clause for technology cells
library unisim ;
use unisim.vcomponents.all;

entity video_buf is 
   port (
      in_data_rsc_z : IN std_logic_vector (2 DOWNTO 0) ;
      in_data_vld_rsc_z : IN std_logic ;
      vga_row_rsc_z : IN std_logic_vector (9 DOWNTO 0) ;
      vga_col_rsc_z : IN std_logic_vector (9 DOWNTO 0) ;
      out_data_rsc_z : OUT std_logic_vector (2 DOWNTO 0) ;
      vga_enable_rsc_z : OUT std_logic ;
      gen_pause_rsc_z : OUT std_logic ;
      clk : IN std_logic ;
      rst : IN std_logic) ;
end video_buf ;

architecture v1 of video_buf is 
   signal buffer_rsc_dualport_addr_1_16, buffer_rsc_dualport_addr_1_15, 
      buffer_rsc_dualport_addr_1_14, buffer_rsc_dualport_addr_1_13, 
      buffer_rsc_dualport_addr_1_12, buffer_rsc_dualport_addr_1_11, nx8332z2, 
      nx48860z1, nx8332z11, nx8332z4, nx8332z12, rd_data2_2, nx7335z2, 
      rd_data2_1, nx6338z2, rd_data2_0: std_logic ;
   
   signal video_buf_core_inst_row_in_sva: std_logic_vector (1 DOWNTO 0) ;
   
   signal video_buf_core_inst_col_in_sva_9, video_buf_core_inst_col_in_sva_8, 
      video_buf_core_inst_col_in_sva_7, video_buf_core_inst_col_in_sva_6, 
      video_buf_core_inst_vga_enable_int_sva_dfm_1, 
      video_buf_core_inst_and_itm_1, nx2364z1, nx2365z1, nx2366z1, nx2367z1, 
      nx2368z1, inc_d_0, nx8474z1, inc_d_1, nx8475z1, inc_d_2, nx8476z1, 
      inc_d_3, nx8477z1, inc_d_4, nx8478z1, inc_d_5, nx8479z1, inc_d_6, 
      nx8480z1, inc_d_7, nx8481z1, inc_d_8, nx51679z1, inc_d_9, 
      video_buf_core_inst_not_row_in_sva_0, nx8539z1, nx8128z1, nx42925z1, 
      nx52268z5, nx8481z2, nx52268z1, nx18093z1, nx8332z5, nx6338z1, 
      nx7335z1, nx8332z3, nx8332z1, nx52268z4, nx52268z3, nx52268z2, 
      nx8332z10, nx8332z9, nx8332z6, nx2368z3, nx2367z3, nx2366z3, nx2365z5, 
      nx2365z4, nx2365z3, nx2364z7, nx2364z6, nx2364z5, nx2364z4, nx2364z3, 
      nx8332z8, nx2363z10, nx2363z9, nx2363z8, nx2363z7, nx2363z6, nx2363z5, 
      nx8332z7, nx2363z4, nx2363z3: std_logic ;
   
   signal DANGLING : std_logic_vector (4 downto 0 );

begin
   modgen_eq_0_eq_muxcy_0 : MUXCY_L port map ( LO=>nx2364z1, CI=>nx8539z1, 
      DI=>nx8481z2, S=>nx2363z3);
   modgen_eq_0_eq_muxcy_1 : MUXCY_L port map ( LO=>nx2365z1, CI=>nx2364z1, 
      DI=>nx8481z2, S=>nx2364z3);
   modgen_eq_0_eq_muxcy_2 : MUXCY_L port map ( LO=>nx2366z1, CI=>nx2365z1, 
      DI=>nx8481z2, S=>nx2365z3);
   modgen_eq_0_eq_muxcy_3 : MUXCY_L port map ( LO=>nx2367z1, CI=>nx2366z1, 
      DI=>nx8481z2, S=>nx2366z3);
   modgen_eq_0_eq_muxcy_4 : MUXCY_L port map ( LO=>nx2368z1, CI=>nx2367z1, 
      DI=>nx8481z2, S=>nx2367z3);
   modgen_eq_0_eq_muxcy_5 : MUXCY port map ( O=>nx8332z11, CI=>nx2368z1, DI
      =>nx8481z2, S=>nx2368z3);
   mem_1 : RAMB16_S4_S4
      generic map (WRITE_MODE_A => "READ_FIRST"
         ,
         WRITE_MODE_B => "WRITE_FIRST") 
       port map ( DOA(3)=>DANGLING(0), DOA(2)=>DANGLING(1), DOA(1)=>DANGLING
      (2), DOA(0)=>DANGLING(3), DOB(3)=>DANGLING(4), DOB(2)=>rd_data2_2, 
      DOB(1)=>rd_data2_1, DOB(0)=>rd_data2_0, ADDRA(11)=>nx8481z2, ADDRA(10)
      =>nx2363z9, ADDRA(9)=>nx2363z4, ADDRA(8)=>nx2364z4, ADDRA(7)=>nx2364z6, 
      ADDRA(6)=>nx2365z4, ADDRA(5)=>buffer_rsc_dualport_addr_1_16, ADDRA(4)
      =>buffer_rsc_dualport_addr_1_15, ADDRA(3)=>
      buffer_rsc_dualport_addr_1_14, ADDRA(2)=>buffer_rsc_dualport_addr_1_13, 
      ADDRA(1)=>buffer_rsc_dualport_addr_1_12, ADDRA(0)=>
      buffer_rsc_dualport_addr_1_11, ADDRB(11)=>nx8481z2, ADDRB(10)=>
      nx2363z6, ADDRB(9)=>nx2363z8, ADDRB(8)=>nx2364z5, ADDRB(7)=>nx2364z7, 
      ADDRB(6)=>nx2365z5, ADDRB(5)=>vga_col_rsc_z(6), ADDRB(4)=>
      vga_col_rsc_z(5), ADDRB(3)=>vga_col_rsc_z(4), ADDRB(2)=>
      vga_col_rsc_z(3), ADDRB(1)=>vga_col_rsc_z(2), ADDRB(0)=>
      vga_col_rsc_z(1), CLKA=>clk, CLKB=>clk, DIA(3)=>nx8481z2, DIA(2)=>
      in_data_rsc_z(2), DIA(1)=>in_data_rsc_z(1), DIA(0)=>in_data_rsc_z(0), 
      DIB(3)=>nx8481z2, DIB(2)=>nx8481z2, DIB(1)=>nx8481z2, DIB(0)=>nx8481z2, 
      ENA=>nx8539z1, ENB=>nx8539z1, SSRA=>nx8481z2, SSRB=>nx8481z2, WEA=>
      nx8332z6, WEB=>nx8481z2);
   reg_q_20 : FDRE port map ( Q=>video_buf_core_inst_col_in_sva_9, C=>clk, 
      CE=>nx18093z1, D=>inc_d_9, R=>nx52268z1);
   reg_q_19 : FDRE port map ( Q=>video_buf_core_inst_col_in_sva_8, C=>clk, 
      CE=>nx18093z1, D=>inc_d_8, R=>nx52268z1);
   reg_q_18 : FDRE port map ( Q=>video_buf_core_inst_col_in_sva_7, C=>clk, 
      CE=>nx18093z1, D=>inc_d_7, R=>nx52268z1);
   reg_q_17 : FDRE port map ( Q=>video_buf_core_inst_col_in_sva_6, C=>clk, 
      CE=>nx18093z1, D=>inc_d_6, R=>nx52268z1);
   reg_q_16 : FDRE port map ( Q=>buffer_rsc_dualport_addr_1_16, C=>clk, CE=>
      nx18093z1, D=>inc_d_5, R=>nx52268z1);
   reg_q_15 : FDRE port map ( Q=>buffer_rsc_dualport_addr_1_15, C=>clk, CE=>
      nx18093z1, D=>inc_d_4, R=>nx52268z1);
   reg_q_14 : FDRE port map ( Q=>buffer_rsc_dualport_addr_1_14, C=>clk, CE=>
      nx18093z1, D=>inc_d_3, R=>nx52268z1);
   reg_q_13 : FDRE port map ( Q=>buffer_rsc_dualport_addr_1_13, C=>clk, CE=>
      nx18093z1, D=>inc_d_2, R=>nx52268z1);
   reg_q_12 : FDRE port map ( Q=>buffer_rsc_dualport_addr_1_12, C=>clk, CE=>
      nx18093z1, D=>inc_d_1, R=>nx52268z1);
   reg_q_11 : FDRE port map ( Q=>buffer_rsc_dualport_addr_1_11, C=>clk, CE=>
      nx18093z1, D=>inc_d_0, R=>nx52268z1);
   xorcy_0 : XORCY port map ( O=>inc_d_0, CI=>nx8539z1, LI=>
      buffer_rsc_dualport_addr_1_11);
   muxcy_0 : MUXCY_L port map ( LO=>nx8474z1, CI=>nx8539z1, DI=>nx8481z2, S
      =>buffer_rsc_dualport_addr_1_11);
   xorcy_1 : XORCY port map ( O=>inc_d_1, CI=>nx8474z1, LI=>
      buffer_rsc_dualport_addr_1_12);
   muxcy_1 : MUXCY_L port map ( LO=>nx8475z1, CI=>nx8474z1, DI=>nx8481z2, S
      =>buffer_rsc_dualport_addr_1_12);
   xorcy_2 : XORCY port map ( O=>inc_d_2, CI=>nx8475z1, LI=>
      buffer_rsc_dualport_addr_1_13);
   muxcy_2 : MUXCY_L port map ( LO=>nx8476z1, CI=>nx8475z1, DI=>nx8481z2, S
      =>buffer_rsc_dualport_addr_1_13);
   xorcy_3 : XORCY port map ( O=>inc_d_3, CI=>nx8476z1, LI=>
      buffer_rsc_dualport_addr_1_14);
   muxcy_3 : MUXCY_L port map ( LO=>nx8477z1, CI=>nx8476z1, DI=>nx8481z2, S
      =>buffer_rsc_dualport_addr_1_14);
   xorcy_4 : XORCY port map ( O=>inc_d_4, CI=>nx8477z1, LI=>
      buffer_rsc_dualport_addr_1_15);
   muxcy_4 : MUXCY_L port map ( LO=>nx8478z1, CI=>nx8477z1, DI=>nx8481z2, S
      =>buffer_rsc_dualport_addr_1_15);
   xorcy_5 : XORCY port map ( O=>inc_d_5, CI=>nx8478z1, LI=>
      buffer_rsc_dualport_addr_1_16);
   muxcy_5 : MUXCY_L port map ( LO=>nx8479z1, CI=>nx8478z1, DI=>nx8481z2, S
      =>buffer_rsc_dualport_addr_1_16);
   xorcy_6 : XORCY port map ( O=>inc_d_6, CI=>nx8479z1, LI=>
      video_buf_core_inst_col_in_sva_6);
   muxcy_6 : MUXCY_L port map ( LO=>nx8480z1, CI=>nx8479z1, DI=>nx8481z2, S
      =>video_buf_core_inst_col_in_sva_6);
   xorcy_7 : XORCY port map ( O=>inc_d_7, CI=>nx8480z1, LI=>
      video_buf_core_inst_col_in_sva_7);
   muxcy_7 : MUXCY_L port map ( LO=>nx8481z1, CI=>nx8480z1, DI=>nx8481z2, S
      =>video_buf_core_inst_col_in_sva_7);
   xorcy_8 : XORCY port map ( O=>inc_d_8, CI=>nx8481z1, LI=>
      video_buf_core_inst_col_in_sva_8);
   muxcy_8 : MUXCY_L port map ( LO=>nx51679z1, CI=>nx8481z1, DI=>nx8481z2, S
      =>video_buf_core_inst_col_in_sva_8);
   xorcy_9 : XORCY port map ( O=>inc_d_9, CI=>nx51679z1, LI=>
      video_buf_core_inst_col_in_sva_9);
   reg_q_1 : FDRE port map ( Q=>video_buf_core_inst_row_in_sva(1), C=>clk, 
      CE=>nx52268z1, D=>nx52268z5, R=>rst);
   reg_q_0 : FDRE port map ( Q=>video_buf_core_inst_row_in_sva(0), C=>clk, 
      CE=>nx52268z1, D=>video_buf_core_inst_not_row_in_sva_0, R=>rst);
   reg_out_data_rsc_mgc_out_stdreg_d_1_2 : FDRE port map ( Q=>
      out_data_rsc_z(2), C=>clk, CE=>nx8332z1, D=>nx8332z3, R=>rst);
   reg_out_data_rsc_mgc_out_stdreg_d_1_1 : FDRE port map ( Q=>
      out_data_rsc_z(1), C=>clk, CE=>nx8332z1, D=>nx7335z1, R=>rst);
   reg_out_data_rsc_mgc_out_stdreg_d_1_0 : FDRE port map ( Q=>
      out_data_rsc_z(0), C=>clk, CE=>nx8332z1, D=>nx6338z1, R=>rst);
   video_buf_core_inst_reg_main_stage_0_2 : FDR port map ( Q=>nx8332z2, C=>
      clk, D=>nx48860z1, R=>rst);
   video_buf_core_inst_reg_vga_enable_int_sva_dfm_1 : FDR port map ( Q=>
      video_buf_core_inst_vga_enable_int_sva_dfm_1, C=>clk, D=>nx42925z1, R
      =>rst);
   video_buf_core_inst_reg_and_itm_1 : FDR port map ( Q=>
      video_buf_core_inst_and_itm_1, C=>clk, D=>nx8128z1, R=>rst);
   video_buf_core_inst_reg_vga_enable_rsc_mgc_out_stdreg_d_drv : FDRE
       port map ( Q=>vga_enable_rsc_z, C=>clk, CE=>nx8332z1, D=>
      video_buf_core_inst_vga_enable_int_sva_dfm_1, R=>rst);
   video_buf_core_inst_reg_gen_pause_rsc_mgc_out_stdreg_d_drv : FDRE
       port map ( Q=>gen_pause_rsc_z, C=>clk, CE=>nx8332z1, D=>
      video_buf_core_inst_and_itm_1, R=>rst);
   video_buf_core_inst_video_buf_core_fsm_inst_reg_state_var : FDR
       port map ( Q=>nx48860z1, C=>clk, D=>nx8539z1, R=>rst);
   ix8332z4325 : FD port map ( Q=>nx8332z4, C=>clk, D=>nx8332z5);
   ix8332z4332 : FD port map ( Q=>nx8332z12, C=>clk, D=>in_data_rsc_z(2));
   ix7335z4324 : FD port map ( Q=>nx7335z2, C=>clk, D=>in_data_rsc_z(1));
   ix6338z4324 : FD port map ( Q=>nx6338z2, C=>clk, D=>in_data_rsc_z(0));
   video_buf_core_inst_not_row_in_sva_0_EXMPLR44 : INV port map ( O=>
      video_buf_core_inst_not_row_in_sva_0, I=>
      video_buf_core_inst_row_in_sva(0));
   ps_vcc : VCC port map ( P=>nx8539z1);
   ix8128z6054 : LUT4
      generic map (INIT => X"1284") 
       port map ( O=>nx8128z1, I0=>vga_row_rsc_z(2), I1=>vga_row_rsc_z(1), 
      I2=>video_buf_core_inst_row_in_sva(1), I3=>
      video_buf_core_inst_row_in_sva(0));
   ix42925z45870 : LUT4
      generic map (INIT => X"AE0C") 
       port map ( O=>nx42925z1, I0=>nx8332z2, I1=>
      video_buf_core_inst_row_in_sva(1), I2=>
      video_buf_core_inst_row_in_sva(0), I3=>
      video_buf_core_inst_vga_enable_int_sva_dfm_1);
   ix52268z1324 : LUT2
      generic map (INIT => X"6") 
       port map ( O=>nx52268z5, I0=>video_buf_core_inst_row_in_sva(1), I1=>
      video_buf_core_inst_row_in_sva(0));
   ps_gnd : GND port map ( G=>nx8481z2);
   ix52268z1186 : LUT4
      generic map (INIT => X"FF80") 
       port map ( O=>nx52268z1, I0=>nx52268z2, I1=>nx52268z3, I2=>nx52268z4, 
      I3=>rst);
   ix18093z1548 : LUT3
      generic map (INIT => X"EA") 
       port map ( O=>nx18093z1, I0=>rst, I1=>in_data_vld_rsc_z, I2=>
      nx48860z1);
   ix8332z1325 : LUT2
      generic map (INIT => X"8") 
       port map ( O=>nx8332z5, I0=>nx8332z6, I1=>nx8332z11);
   ix6338z1530 : LUT3
      generic map (INIT => X"D8") 
       port map ( O=>nx6338z1, I0=>nx8332z4, I1=>nx6338z2, I2=>rd_data2_0);
   ix7335z1530 : LUT3
      generic map (INIT => X"D8") 
       port map ( O=>nx7335z1, I0=>nx8332z4, I1=>nx7335z2, I2=>rd_data2_1);
   ix8332z1531 : LUT3
      generic map (INIT => X"D8") 
       port map ( O=>nx8332z3, I0=>nx8332z4, I1=>nx8332z12, I2=>rd_data2_2);
   ix8332z1322 : LUT2
      generic map (INIT => X"8") 
       port map ( O=>nx8332z1, I0=>nx8332z2, I1=>nx48860z1);
   ix52268z1445 : LUT4
      generic map (INIT => X"0080") 
       port map ( O=>nx52268z4, I0=>in_data_vld_rsc_z, I1=>
      buffer_rsc_dualport_addr_1_13, I2=>nx48860z1, I3=>
      video_buf_core_inst_col_in_sva_6);
   ix52268z34084 : LUT4
      generic map (INIT => X"8000") 
       port map ( O=>nx52268z3, I0=>buffer_rsc_dualport_addr_1_16, I1=>
      buffer_rsc_dualport_addr_1_15, I2=>buffer_rsc_dualport_addr_1_14, I3=>
      buffer_rsc_dualport_addr_1_12);
   ix52268z1347 : LUT4
      generic map (INIT => X"0020") 
       port map ( O=>nx52268z2, I0=>buffer_rsc_dualport_addr_1_11, I1=>
      video_buf_core_inst_col_in_sva_9, I2=>video_buf_core_inst_col_in_sva_8, 
      I3=>video_buf_core_inst_col_in_sva_7);
   ix8332z1330 : LUT2
      generic map (INIT => X"8") 
       port map ( O=>nx8332z10, I0=>in_data_vld_rsc_z, I1=>nx48860z1);
   ix8332z42409 : LUT4
      generic map (INIT => X"A080") 
       port map ( O=>nx8332z9, I0=>video_buf_core_inst_row_in_sva(1), I1=>
      video_buf_core_inst_row_in_sva(0), I2=>
      video_buf_core_inst_col_in_sva_9, I3=>video_buf_core_inst_col_in_sva_8
   );
   ix8332z8230 : LUT4
      generic map (INIT => X"1B00") 
       port map ( O=>nx8332z6, I0=>nx8332z7, I1=>nx8332z8, I2=>nx8332z9, I3
      =>nx8332z10);
   ix2368z1324 : LUT2
      generic map (INIT => X"9") 
       port map ( O=>nx2368z3, I0=>buffer_rsc_dualport_addr_1_11, I1=>
      vga_col_rsc_z(1));
   ix2367z35140 : LUT4
      generic map (INIT => X"8421") 
       port map ( O=>nx2367z3, I0=>buffer_rsc_dualport_addr_1_13, I1=>
      buffer_rsc_dualport_addr_1_12, I2=>vga_col_rsc_z(3), I3=>
      vga_col_rsc_z(2));
   ix2366z35140 : LUT4
      generic map (INIT => X"8421") 
       port map ( O=>nx2366z3, I0=>buffer_rsc_dualport_addr_1_15, I1=>
      buffer_rsc_dualport_addr_1_14, I2=>vga_col_rsc_z(5), I3=>
      vga_col_rsc_z(4));
   ix2365z1323 : LUT2
      generic map (INIT => X"6") 
       port map ( O=>nx2365z5, I0=>vga_row_rsc_z(1), I1=>vga_col_rsc_z(7));
   ix2365z1322 : LUT2
      generic map (INIT => X"6") 
       port map ( O=>nx2365z4, I0=>video_buf_core_inst_row_in_sva(0), I1=>
      video_buf_core_inst_col_in_sva_6);
   ix2365z38188 : LUT4
      generic map (INIT => X"9009") 
       port map ( O=>nx2365z3, I0=>nx2365z4, I1=>nx2365z5, I2=>
      buffer_rsc_dualport_addr_1_16, I3=>vga_col_rsc_z(6));
   ix2364z39809 : LUT4
      generic map (INIT => X"965A") 
       port map ( O=>nx2364z7, I0=>vga_row_rsc_z(2), I1=>vga_row_rsc_z(1), 
      I2=>vga_col_rsc_z(8), I3=>vga_col_rsc_z(7));
   ix2364z39808 : LUT4
      generic map (INIT => X"965A") 
       port map ( O=>nx2364z6, I0=>video_buf_core_inst_row_in_sva(1), I1=>
      video_buf_core_inst_row_in_sva(0), I2=>
      video_buf_core_inst_col_in_sva_7, I3=>video_buf_core_inst_col_in_sva_6
   );
   ix2364z1422 : LUT3
      generic map (INIT => X"69") 
       port map ( O=>nx2364z5, I0=>nx2363z7, I1=>vga_row_rsc_z(1), I2=>
      vga_col_rsc_z(9));
   ix2364z1421 : LUT3
      generic map (INIT => X"69") 
       port map ( O=>nx2364z4, I0=>nx8332z7, I1=>
      video_buf_core_inst_row_in_sva(0), I2=>
      video_buf_core_inst_col_in_sva_8);
   ix2364z38188 : LUT4
      generic map (INIT => X"9009") 
       port map ( O=>nx2364z3, I0=>nx2364z4, I1=>nx2364z5, I2=>nx2364z6, I3
      =>nx2364z7);
   ix8332z60872 : LUT4
      generic map (INIT => X"E8A0") 
       port map ( O=>nx8332z8, I0=>video_buf_core_inst_row_in_sva(1), I1=>
      video_buf_core_inst_row_in_sva(0), I2=>
      video_buf_core_inst_col_in_sva_9, I3=>video_buf_core_inst_col_in_sva_8
   );
   ix2363z19 : LUT4
      generic map (INIT => X"FAE8") 
       port map ( O=>nx2363z10, I0=>video_buf_core_inst_row_in_sva(1), I1=>
      video_buf_core_inst_row_in_sva(0), I2=>
      video_buf_core_inst_col_in_sva_9, I3=>video_buf_core_inst_col_in_sva_8
   );
   ix2363z1550 : LUT3
      generic map (INIT => X"E4") 
       port map ( O=>nx2363z9, I0=>nx8332z7, I1=>nx2363z10, I2=>nx8332z8);
   ix2363z16069 : LUT4
      generic map (INIT => X"399C") 
       port map ( O=>nx2363z8, I0=>nx2363z7, I1=>vga_row_rsc_z(2), I2=>
      vga_row_rsc_z(1), I3=>vga_col_rsc_z(9));
   ix2363z7303 : LUT4
      generic map (INIT => X"175F") 
       port map ( O=>nx2363z7, I0=>vga_row_rsc_z(2), I1=>vga_row_rsc_z(1), 
      I2=>vga_col_rsc_z(8), I3=>vga_col_rsc_z(7));
   ix2363z51559 : LUT4
      generic map (INIT => X"C440") 
       port map ( O=>nx2363z6, I0=>nx2363z7, I1=>vga_row_rsc_z(2), I2=>
      vga_row_rsc_z(1), I3=>vga_col_rsc_z(9));
   ix2363z1324 : LUT2
      generic map (INIT => X"6") 
       port map ( O=>nx2363z5, I0=>video_buf_core_inst_row_in_sva(1), I1=>
      video_buf_core_inst_col_in_sva_9);
   ix8332z7302 : LUT4
      generic map (INIT => X"175F") 
       port map ( O=>nx8332z7, I0=>video_buf_core_inst_row_in_sva(1), I1=>
      video_buf_core_inst_row_in_sva(0), I2=>
      video_buf_core_inst_col_in_sva_7, I3=>video_buf_core_inst_col_in_sva_6
   );
   ix2363z16065 : LUT4
      generic map (INIT => X"399C") 
       port map ( O=>nx2363z4, I0=>nx8332z7, I1=>nx2363z5, I2=>
      video_buf_core_inst_row_in_sva(0), I3=>
      video_buf_core_inst_col_in_sva_8);
   ix2363z35141 : LUT4
      generic map (INIT => X"8421") 
       port map ( O=>nx2363z3, I0=>nx2363z4, I1=>nx2363z6, I2=>nx2363z8, I3
      =>nx2363z9);
end v1 ;

